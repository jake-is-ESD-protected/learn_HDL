/*
*****************************************************************************************
project name:       dreg
auth:               Jakob Tschavoll
date:               03.11.21
brief:              system verilog testbench for D-FF
version:            V1.0
*****************************************************************************************
*/