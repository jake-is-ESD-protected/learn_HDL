/*
*****************************************************************************************
project name:       ram16k_verilog
auth:               Jakob Tschavoll
date:               03.11.21
brief:              system verilog testbench for RAM
version:            V1.0
*****************************************************************************************
*/