/*
*****************************************************************************************
project name:       pcount
auth:               Jakob Tschavoll
date:               03.11.21
brief:              system verilog implementation of a counter
version:            V1.0
*****************************************************************************************
*/