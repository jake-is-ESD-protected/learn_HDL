/*
*****************************************************************************************
project name:       pcount
auth:               Jakob Tschavoll
date:               03.11.21
brief:              system verilog testbench for counter
version:            V1.0
*****************************************************************************************
*/